// when controling mux_ui module, after each ui, a clear must be called before the 
// next change_instruction goes high;
// each clear must be called high after done is high

module process_game ();


endmodule // process_game




